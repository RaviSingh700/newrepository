module tb;
endmodule
